interface jtag_if;
    logic trst_n;
    logic tck;
    logic tms;
    logic tdi;
    logic tdo;
    logic tdo_en;
endinterface //jtag_if