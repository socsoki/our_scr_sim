//-----------------------------------------------------------------
//                     Basic Peripheral SoC
//                           V1.1
//                     Ultra-Embedded.com
//                     Copyright 2014-2020
//
//                 Email: admin@ultra-embedded.com
//
//                         License: GPL
// If you would like a version with a more permissive license for
// use in closed source commercial applications please contact me
// for details.
//-----------------------------------------------------------------
//
// This file is open source HDL; you can redistribute it and/or 
// modify it under the terms of the GNU General Public License as 
// published by the Free Software Foundation; either version 2 of 
// the License, or (at your option) any later version.
//
// This file is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public 
// License along with this file; if not, write to the Free Software
// Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA 02111-1307
// USA
//-----------------------------------------------------------------

//-----------------------------------------------------------------
//                          Generated File
//-----------------------------------------------------------------

`define ULITE_RX    8'h0

    `define ULITE_RX_DATA_DEFAULT    0
    `define ULITE_RX_DATA_B          0
    `define ULITE_RX_DATA_T          7
    `define ULITE_RX_DATA_W          8
    `define ULITE_RX_DATA_R          7:0

`define ULITE_TX    8'h4

    `define ULITE_TX_DATA_DEFAULT    0
    `define ULITE_TX_DATA_B          0
    `define ULITE_TX_DATA_T          7
    `define ULITE_TX_DATA_W          8
    `define ULITE_TX_DATA_R          7:0

`define ULITE_STATUS    8'h8

    `define ULITE_STATUS_IE      4
    `define ULITE_STATUS_IE_DEFAULT    0
    `define ULITE_STATUS_IE_B          4
    `define ULITE_STATUS_IE_T          4
    `define ULITE_STATUS_IE_W          1
    `define ULITE_STATUS_IE_R          4:4

    `define ULITE_STATUS_TXFULL      3
    `define ULITE_STATUS_TXFULL_DEFAULT    0
    `define ULITE_STATUS_TXFULL_B          3
    `define ULITE_STATUS_TXFULL_T          3
    `define ULITE_STATUS_TXFULL_W          1
    `define ULITE_STATUS_TXFULL_R          3:3

    `define ULITE_STATUS_TXEMPTY      2
    `define ULITE_STATUS_TXEMPTY_DEFAULT    0
    `define ULITE_STATUS_TXEMPTY_B          2
    `define ULITE_STATUS_TXEMPTY_T          2
    `define ULITE_STATUS_TXEMPTY_W          1
    `define ULITE_STATUS_TXEMPTY_R          2:2

    `define ULITE_STATUS_RXFULL      1
    `define ULITE_STATUS_RXFULL_DEFAULT    0
    `define ULITE_STATUS_RXFULL_B          1
    `define ULITE_STATUS_RXFULL_T          1
    `define ULITE_STATUS_RXFULL_W          1
    `define ULITE_STATUS_RXFULL_R          1:1

    `define ULITE_STATUS_RXVALID      0
    `define ULITE_STATUS_RXVALID_DEFAULT    0
    `define ULITE_STATUS_RXVALID_B          0
    `define ULITE_STATUS_RXVALID_T          0
    `define ULITE_STATUS_RXVALID_W          1
    `define ULITE_STATUS_RXVALID_R          0:0

`define ULITE_CONTROL    8'hc

    `define ULITE_CONTROL_IE      4
    `define ULITE_CONTROL_IE_DEFAULT    0
    `define ULITE_CONTROL_IE_B          4
    `define ULITE_CONTROL_IE_T          4
    `define ULITE_CONTROL_IE_W          1
    `define ULITE_CONTROL_IE_R          4:4

    `define ULITE_CONTROL_RST_RX      1
    `define ULITE_CONTROL_RST_RX_DEFAULT    0
    `define ULITE_CONTROL_RST_RX_B          1
    `define ULITE_CONTROL_RST_RX_T          1
    `define ULITE_CONTROL_RST_RX_W          1
    `define ULITE_CONTROL_RST_RX_R          1:1

    `define ULITE_CONTROL_RST_TX      0
    `define ULITE_CONTROL_RST_TX_DEFAULT    0
    `define ULITE_CONTROL_RST_TX_B          0
    `define ULITE_CONTROL_RST_TX_T          0
    `define ULITE_CONTROL_RST_TX_W          1
    `define ULITE_CONTROL_RST_TX_R          0:0

//-----------------------------------------------------------------
// Module:  UART (uartlite compatable)
//-----------------------------------------------------------------
module uart_lite
//-----------------------------------------------------------------
// Params
//-----------------------------------------------------------------
#(
     parameter CLK_FREQ         = 1843200
    ,parameter BAUDRATE         = 115200
)
//-----------------------------------------------------------------
// Ports
//-----------------------------------------------------------------
(
    // Inputs
     input          clk_i
    ,input          rst_i
    ,input          cfg_awvalid_i
    ,input  [31:0]  cfg_awaddr_i
    ,input          cfg_wvalid_i
    ,input  [31:0]  cfg_wdata_i
    ,input  [3:0]   cfg_wstrb_i
    ,input          cfg_bready_i
    ,input          cfg_arvalid_i
    ,input  [31:0]  cfg_araddr_i
    ,input          cfg_rready_i
    ,input          rx_i

    // Outputs
    ,output         cfg_awready_o
    ,output         cfg_wready_o
    ,output         cfg_bvalid_o
    ,output [1:0]   cfg_bresp_o
    ,output         cfg_arready_o
    ,output         cfg_rvalid_o
    ,output [31:0]  cfg_rdata_o
    ,output [1:0]   cfg_rresp_o
    ,output         tx_o
    ,output         intr_o
);

//-----------------------------------------------------------------
// Write address / data split
//-----------------------------------------------------------------
// Address but no data ready
reg awvalid_q;

// Data but no data ready
reg wvalid_q;

wire wr_cmd_accepted_w  = (cfg_awvalid_i && cfg_awready_o) || awvalid_q;
wire wr_data_accepted_w = (cfg_wvalid_i  && cfg_wready_o)  || wvalid_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    awvalid_q <= 1'b0;
else if (cfg_awvalid_i && cfg_awready_o && !wr_data_accepted_w)
    awvalid_q <= 1'b1;
else if (wr_data_accepted_w)
    awvalid_q <= 1'b0;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    wvalid_q <= 1'b0;
else if (cfg_wvalid_i && cfg_wready_o && !wr_cmd_accepted_w)
    wvalid_q <= 1'b1;
else if (wr_cmd_accepted_w)
    wvalid_q <= 1'b0;

//-----------------------------------------------------------------
// Capture address (for delayed data)
//-----------------------------------------------------------------
reg [7:0] wr_addr_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    wr_addr_q <= 8'b0;
else if (cfg_awvalid_i && cfg_awready_o)
    wr_addr_q <= cfg_awaddr_i[7:0];

wire [7:0] wr_addr_w = awvalid_q ? wr_addr_q : cfg_awaddr_i[7:0];

//-----------------------------------------------------------------
// Retime write data
//-----------------------------------------------------------------
reg [31:0] wr_data_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    wr_data_q <= 32'b0;
else if (cfg_wvalid_i && cfg_wready_o)
    wr_data_q <= cfg_wdata_i;

//-----------------------------------------------------------------
// Request Logic
//-----------------------------------------------------------------
wire read_en_w  = cfg_arvalid_i & cfg_arready_o;
wire write_en_w = wr_cmd_accepted_w && wr_data_accepted_w;

//-----------------------------------------------------------------
// Accept Logic
//-----------------------------------------------------------------
assign cfg_arready_o = ~cfg_rvalid_o;
assign cfg_awready_o = ~cfg_bvalid_o && ~cfg_arvalid_i && ~awvalid_q;
assign cfg_wready_o  = ~cfg_bvalid_o && ~cfg_arvalid_i && ~wvalid_q;


//-----------------------------------------------------------------
// Register ulite_rx
//-----------------------------------------------------------------
reg ulite_rx_wr_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_rx_wr_q <= 1'b0;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_RX))
    ulite_rx_wr_q <= 1'b1;
else
    ulite_rx_wr_q <= 1'b0;


//-----------------------------------------------------------------
// Register ulite_tx
//-----------------------------------------------------------------
reg ulite_tx_wr_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_tx_wr_q <= 1'b0;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_TX))
    ulite_tx_wr_q <= 1'b1;
else
    ulite_tx_wr_q <= 1'b0;

// ulite_tx_data [external]
wire [7:0]  ulite_tx_data_out_w = wr_data_q[`ULITE_TX_DATA_R];


//-----------------------------------------------------------------
// Register ulite_status
//-----------------------------------------------------------------
reg ulite_status_wr_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_status_wr_q <= 1'b0;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_STATUS))
    ulite_status_wr_q <= 1'b1;
else
    ulite_status_wr_q <= 1'b0;

//-----------------------------------------------------------------
// Register ulite_control
//-----------------------------------------------------------------
reg ulite_control_wr_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_control_wr_q <= 1'b0;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_CONTROL))
    ulite_control_wr_q <= 1'b1;
else
    ulite_control_wr_q <= 1'b0;

// ulite_control_ie [internal]
reg        ulite_control_ie_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_control_ie_q <= 1'd`ULITE_CONTROL_IE_DEFAULT;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_CONTROL))
    ulite_control_ie_q <= cfg_wdata_i[`ULITE_CONTROL_IE_R];

wire        ulite_control_ie_out_w = ulite_control_ie_q;


// ulite_control_rst_rx [auto_clr]
reg        ulite_control_rst_rx_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_control_rst_rx_q <= 1'd`ULITE_CONTROL_RST_RX_DEFAULT;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_CONTROL))
    ulite_control_rst_rx_q <= cfg_wdata_i[`ULITE_CONTROL_RST_RX_R];
else
    ulite_control_rst_rx_q <= 1'd`ULITE_CONTROL_RST_RX_DEFAULT;

wire        ulite_control_rst_rx_out_w = ulite_control_rst_rx_q;


// ulite_control_rst_tx [auto_clr]
reg        ulite_control_rst_tx_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    ulite_control_rst_tx_q <= 1'd`ULITE_CONTROL_RST_TX_DEFAULT;
else if (write_en_w && (wr_addr_w[7:0] == `ULITE_CONTROL))
    ulite_control_rst_tx_q <= cfg_wdata_i[`ULITE_CONTROL_RST_TX_R];
else
    ulite_control_rst_tx_q <= 1'd`ULITE_CONTROL_RST_TX_DEFAULT;

wire        ulite_control_rst_tx_out_w = ulite_control_rst_tx_q;


wire [7:0]  ulite_rx_data_in_w;
wire        ulite_status_ie_in_w;
wire        ulite_status_txfull_in_w;
wire        ulite_status_txempty_in_w;
wire        ulite_status_rxfull_in_w;
wire        ulite_status_rxvalid_in_w;


//-----------------------------------------------------------------
// Read mux
//-----------------------------------------------------------------
reg [31:0] data_r;

always @ *
begin
    data_r = 32'b0;

    case (cfg_araddr_i[7:0])

    `ULITE_RX:
    begin
        data_r[`ULITE_RX_DATA_R] = ulite_rx_data_in_w;
    end
    `ULITE_STATUS:
    begin
        data_r[`ULITE_STATUS_IE_R] = ulite_status_ie_in_w;
        data_r[`ULITE_STATUS_TXFULL_R] = ulite_status_txfull_in_w;
        data_r[`ULITE_STATUS_TXEMPTY_R] = ulite_status_txempty_in_w;
        data_r[`ULITE_STATUS_RXFULL_R] = ulite_status_rxfull_in_w;
        data_r[`ULITE_STATUS_RXVALID_R] = ulite_status_rxvalid_in_w;
    end
    `ULITE_CONTROL:
    begin
        data_r[`ULITE_CONTROL_IE_R] = ulite_control_ie_q;
    end
    default :
        data_r = 32'b0;
    endcase
end

//-----------------------------------------------------------------
// RVALID
//-----------------------------------------------------------------
reg rvalid_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    rvalid_q <= 1'b0;
else if (read_en_w)
    rvalid_q <= 1'b1;
else if (cfg_rready_i)
    rvalid_q <= 1'b0;

assign cfg_rvalid_o = rvalid_q;

//-----------------------------------------------------------------
// Retime read response
//-----------------------------------------------------------------
reg [31:0] rd_data_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    rd_data_q <= 32'b0;
else if (!cfg_rvalid_o || cfg_rready_i)
    rd_data_q <= data_r;

assign cfg_rdata_o = rd_data_q;
assign cfg_rresp_o = 2'b0;

//-----------------------------------------------------------------
// BVALID
//-----------------------------------------------------------------
reg bvalid_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    bvalid_q <= 1'b0;
else if (write_en_w)
    bvalid_q <= 1'b1;
else if (cfg_bready_i)
    bvalid_q <= 1'b0;

assign cfg_bvalid_o = bvalid_q;
assign cfg_bresp_o  = 2'b0;

wire ulite_rx_rd_req_w = read_en_w & (cfg_araddr_i[7:0] == `ULITE_RX);

wire ulite_rx_wr_req_w = ulite_rx_wr_q;
wire ulite_tx_wr_req_w = ulite_tx_wr_q;

//-----------------------------------------------------------------
// Registers
//-----------------------------------------------------------------

// Configuration
localparam   STOP_BITS = 1'b0; // 0 = 1, 1 = 2
localparam   BIT_DIV   = (CLK_FREQ / BAUDRATE) - 1;

localparam   START_BIT = 4'd0;
localparam   STOP_BIT0 = 4'd9;
localparam   STOP_BIT1 = 4'd10;

// Xilinx placement pragmas:
//synthesis attribute IOB of txd_q is "TRUE"

// TX Signals
reg          tx_busy_q;
reg [3:0]    tx_bits_q;
reg [31:0]   tx_count_q;
reg [7:0]    tx_shift_reg_q;
reg          txd_q;

// RX Signals
reg          rxd_q;
reg [7:0]    rx_data_q;
reg [3:0]    rx_bits_q;
reg [31:0]   rx_count_q;
reg [7:0]    rx_shift_reg_q;
reg          rx_ready_q;
reg          rx_busy_q;

reg          rx_err_q;

//-----------------------------------------------------------------
// Re-sync RXD
//-----------------------------------------------------------------
reg rxd_ms_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
begin
   rxd_ms_q <= 1'b1;
   rxd_q    <= 1'b1;
end
else
begin
   rxd_ms_q <= rx_i;
   rxd_q    <= rxd_ms_q;
end

//-----------------------------------------------------------------
// RX Clock Divider
//-----------------------------------------------------------------
wire rx_sample_w = (rx_count_q == 32'b0);

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    rx_count_q        <= 32'b0;
else
begin
    // Inactive
    if (!rx_busy_q)
        rx_count_q    <= {1'b0, BIT_DIV[31:1]};
    // Rx bit timer
    else if (rx_count_q != 0)
        rx_count_q    <= (rx_count_q - 1);
    // Active
    else if (rx_sample_w)
    begin
        // Last bit?
        if ((rx_bits_q == STOP_BIT0 && !STOP_BITS) || (rx_bits_q == STOP_BIT1 && STOP_BITS))
            rx_count_q    <= 32'b0;
        else
            rx_count_q    <= BIT_DIV;
    end
end

//-----------------------------------------------------------------
// RX Shift Register
//-----------------------------------------------------------------
always @ (posedge clk_i or posedge rst_i)
if (rst_i)
begin
    rx_shift_reg_q <= 8'h00;
    rx_busy_q      <= 1'b0;
end
// Rx busy
else if (rx_busy_q && rx_sample_w)
begin
    // Last bit?
    if (rx_bits_q == STOP_BIT0 && !STOP_BITS)
        rx_busy_q <= 1'b0;
    else if (rx_bits_q == STOP_BIT1 && STOP_BITS)
        rx_busy_q <= 1'b0;
    else if (rx_bits_q == START_BIT)
    begin
        // Start bit should still be low as sampling mid
        // way through start bit, so if high, error!
        if (rxd_q)
            rx_busy_q <= 1'b0;
    end
    // Rx shift register
    else 
        rx_shift_reg_q <= {rxd_q, rx_shift_reg_q[7:1]};
end
// Start bit?
else if (!rx_busy_q && rxd_q == 1'b0)
begin
    rx_shift_reg_q <= 8'h00;
    rx_busy_q      <= 1'b1;
end

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    rx_bits_q  <= START_BIT;
else if (rx_sample_w && rx_busy_q)
begin
    if ((rx_bits_q == STOP_BIT1 && STOP_BITS) || (rx_bits_q == STOP_BIT0 && !STOP_BITS))
        rx_bits_q <= START_BIT;
    else
        rx_bits_q <= rx_bits_q + 4'd1;
end
else if (!rx_busy_q && (BIT_DIV == 32'b0))
    rx_bits_q  <= START_BIT + 4'd1;
else if (!rx_busy_q)
    rx_bits_q  <= START_BIT;

//-----------------------------------------------------------------
// RX Data
//-----------------------------------------------------------------
always @ (posedge clk_i or posedge rst_i)
if (rst_i)
begin
   rx_ready_q      <= 1'b0;
   rx_data_q       <= 8'h00;
   rx_err_q        <= 1'b0;
end
else
begin
   // If reading data, reset data state
   if (ulite_rx_rd_req_w || ulite_control_rst_rx_out_w)
   begin
       rx_ready_q <= 1'b0;
       rx_err_q   <= 1'b0;
   end

   if (rx_busy_q && rx_sample_w)
   begin
       // Stop bit
       if ((rx_bits_q == STOP_BIT1 && STOP_BITS) || (rx_bits_q == STOP_BIT0 && !STOP_BITS))
       begin
           // RXD should be still high
           if (rxd_q)
           begin
               rx_data_q      <= rx_shift_reg_q;
               rx_ready_q     <= 1'b1;
           end
           // Bad Stop bit - wait for a full bit period
           // before allowing start bit detection again
           else
           begin
               rx_ready_q      <= 1'b0;
               rx_data_q       <= 8'h00;
               rx_err_q        <= 1'b1;
           end
       end
       // Mid start bit sample - if high then error
       else if (rx_bits_q == START_BIT && rxd_q)
           rx_err_q        <= 1'b1;
   end
end

assign ulite_rx_data_in_w        = rx_data_q;
assign ulite_status_rxvalid_in_w = rx_ready_q;
assign ulite_status_rxfull_in_w  = rx_ready_q;

//-----------------------------------------------------------------
// TX Clock Divider
//-----------------------------------------------------------------
wire tx_sample_w = (tx_count_q == 32'b0);

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    tx_count_q      <= 32'b0;
else
begin
    // Idle
    if (!tx_busy_q)
        tx_count_q  <= BIT_DIV;
    // Tx bit timer
    else if (tx_count_q != 0)
        tx_count_q  <= (tx_count_q - 1);
    else if (tx_sample_w)
        tx_count_q  <= BIT_DIV;
end

//-----------------------------------------------------------------
// TX Shift Register
//-----------------------------------------------------------------
reg tx_complete_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
begin
    tx_shift_reg_q <= 8'h00;
    tx_busy_q      <= 1'b0;
    tx_complete_q  <= 1'b0;
end
// Tx busy
else if (tx_busy_q)
begin
    // Shift tx data
    if (tx_bits_q != START_BIT && tx_sample_w)
        tx_shift_reg_q <= {1'b0, tx_shift_reg_q[7:1]};

    // Last bit?
    if (tx_bits_q == STOP_BIT0 && tx_sample_w && !STOP_BITS)
    begin
        tx_busy_q      <= 1'b0;
        tx_complete_q  <= 1'b1;
    end
    else if (tx_bits_q == STOP_BIT1 && tx_sample_w && STOP_BITS)
    begin
        tx_busy_q      <= 1'b0;
        tx_complete_q  <= 1'b1;
    end
end
// Buffer data to transmit
else if (ulite_tx_wr_req_w)
begin
    tx_shift_reg_q <= ulite_tx_data_out_w;
    tx_busy_q      <= 1'b1;
    tx_complete_q  <= 1'b0;
end
else
    tx_complete_q  <= 1'b0;

assign ulite_status_txfull_in_w  = tx_busy_q;
assign ulite_status_txempty_in_w = ~tx_busy_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    tx_bits_q  <= 4'd0;
else if (tx_sample_w && tx_busy_q)
begin
    if ((tx_bits_q == STOP_BIT1 && STOP_BITS) || (tx_bits_q == STOP_BIT0 && !STOP_BITS))
        tx_bits_q <= START_BIT;
    else
        tx_bits_q <= tx_bits_q + 4'd1;
end

//-----------------------------------------------------------------
// UART Tx Pin
//-----------------------------------------------------------------
reg txd_r;

always @ *
begin
    txd_r = 1'b1;

    if (tx_busy_q)
    begin
        // Start bit (TXD = L)
        if (tx_bits_q == START_BIT)
            txd_r = 1'b0;
        // Stop bits (TXD = H)
        else if (tx_bits_q == STOP_BIT0 || tx_bits_q == STOP_BIT1)
            txd_r = 1'b1;
        // Data bits
        else
            txd_r = tx_shift_reg_q[0];
    end
end

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
    txd_q <= 1'b1;
else
    txd_q <= txd_r;

assign tx_o = txd_q;

//-----------------------------------------------------------------
// Interrupt
//-----------------------------------------------------------------
reg intr_q;

always @ (posedge clk_i or posedge rst_i)
if (rst_i)
   intr_q <= 1'b0;
else if (tx_complete_q)
   intr_q <= 1'b1;
else if (ulite_status_rxvalid_in_w)
   intr_q <= 1'b1;
else
   intr_q <= 1'b0;

assign ulite_status_ie_in_w = ulite_control_ie_out_w;

//-----------------------------------------------------------------
// Assignments
//-----------------------------------------------------------------
assign intr_o = intr_q;


endmodule